`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: CSULB
// Engineers: Jose Aceves & Amin Rezaei 
// Create Date: 11/09/2020 10:16:17 PM
// Design Name: 361_Lab5
// Module Name: Circuit_SA1
//////////////////////////////////////////////////////////////////////////////////

module Circuit_SA1(
    input A,
    input B,
    input C,
    output F0,
    output F1
    );
        
    wire F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBllANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep;
    wire F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep;
    wire F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k11bTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep;
    wire F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz11WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep;
    wire F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehlUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep;
    wire F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwlD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep;
    wire F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph115BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep;
    wire F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1blTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep;
    
    assign F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBllANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep = A;
    assign F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep = B;
    assign F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k11bTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep = C;
    assign F0=F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz11WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep;
    assign F1=F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehlUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep;
    assign F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwlD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep=F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBllANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep^F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep;
    assign F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz11WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep=F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwlD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep^F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k11bTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep;
    assign F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph115BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep=F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k11bTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep&(F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwlD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep|~F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwlD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep);      
    assign F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1blTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep=F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBllANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep&F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep;
    assign F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehlUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep=F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1bTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph115BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep|F1eC$svu81nh5pK4dITXDZZsuEujVZQxJv8gL2H$Z_DVeR0hZrD5waPcOhCBxrmeuY1TiPwLaN3FpVmIeJMjyBHiqDgavei0A1GmpKAHZEw_FQn_PFmMdOBa_HgFlDE0PDuKId5HRfKJfnGI4pCdcv0Ix0KL$$_lzIr5J4n9gx5UdDBL24WftmjCC8A$t3fznDO4al_n5ycKxxpHC_dsl6sEmO2BIyRqgBMkgOTXli5E0VdPr23SGiFREvJepR1xuPIntruwO12Xvj50CNj8q4$BC5EwPx7TgmIzv3qwJ8LWeV6hRAEA$H8WXjnlfz1WEGE45aeIO6eiRDRe5WQVy3qDdS5LaMZqI4vT6ZR7dgF1gestwehUoaQkl3aeGofG6HkSIg5$iKT6jRv31YNuGrad1t6k1blTpE81TyLrKdWbBlANEwpGIwD3kGQyQ6YNserEMvosR6Ph15BzCfIbRJqAlmHgPjqaGyYFUmMxqVjXaysEyCmNstmvsRil2GXep;
      
endmodule
